-- Se implementa un flip flop de tipo RS